-- Librerie utilizzate
library IEEE;
use IEEE.std_logic_1164.all;
entity testbench_new is
end testbench_new;
-- Dichiarazione dell'entit�
architecture interleaver_test of testbench_new is
	component interleaver
   generic(Nbit: POSITIVE := 1024);
		port (
			clock		: in std_logic;						-- segnale di clock
			reset	: in std_logic;							-- segnale di reset
			bit_in		: in std_logic;	-- ingresso
			bit_out 	: out std_logic	-- uscita
			);
	end component;
-----------------------------------------------------
--CONSTANT
	CONSTANT clock_period : TIME := 8 ns;
	CONSTANT len : INTEGER := 2050;
	--INPUT SIGNALS
	SIGNAL clock_tb : std_logic := '0';
	SIGNAL reset_tb : std_logic := '1';
	SIGNAL bit_in_tb : std_logic := '0';


	--OUTPUT SIGNALS2
	SIGNAL bit_out_tb : std_logic := '0';

	SIGNAL testing: Boolean :=True;

	signal count: INTEGER:= 0;

	BEGIN
		I: interleaver
       generic map(Nbit => 1024)
       PORT MAP
           (clock => clock_tb, reset => reset_tb, bit_in => bit_in_tb, bit_out =>bit_out_tb);

--Generates clk
	clock_tb <=NOT clock_tb AFTER clock_period/2 WHEN testing ELSE '0';
    reset_tb <= '0' after 2*clock_Period;

    --Runs simulation for len cycles
    proc_test: process(clock_tb, reset_tb)

    begin

        if(reset_tb = '1') then
				bit_in_tb <= '0';
               count <= -1;

       elsif rising_edge(clock_tb) then
           CASE count IS
                WHEN 0 => bit_in_tb <= '1';
                WHEN 1 => bit_in_tb <= '1';
                WHEN 2 => bit_in_tb <= '1';
                WHEN 3 => bit_in_tb <= '1';
                WHEN 4 => bit_in_tb <= '1';
                WHEN 5 => bit_in_tb <= '1';
                WHEN 6 => bit_in_tb <= '0';
                WHEN 7 => bit_in_tb <= '1';
                WHEN 8 => bit_in_tb <= '0';
                WHEN 9 => bit_in_tb <= '0';
                WHEN 10 => bit_in_tb <= '1';
                WHEN 11 => bit_in_tb <= '1';
                WHEN 12 => bit_in_tb <= '0';
                WHEN 13 => bit_in_tb <= '0';
                WHEN 14 => bit_in_tb <= '1';
                WHEN 15 => bit_in_tb <= '1';
                WHEN 16 => bit_in_tb <= '0';
                WHEN 17 => bit_in_tb <= '1';
                WHEN 18 => bit_in_tb <= '1';
                WHEN 19 => bit_in_tb <= '1';
                WHEN 20 => bit_in_tb <= '0';
                WHEN 21 => bit_in_tb <= '0';
                WHEN 22 => bit_in_tb <= '0';
                WHEN 23 => bit_in_tb <= '0';
                WHEN 24 => bit_in_tb <= '1';
                WHEN 25 => bit_in_tb <= '0';
                WHEN 26 => bit_in_tb <= '0';
                WHEN 27 => bit_in_tb <= '1';
                WHEN 28 => bit_in_tb <= '0';
                WHEN 29 => bit_in_tb <= '1';
                WHEN 30 => bit_in_tb <= '0';
                WHEN 31 => bit_in_tb <= '1';
                WHEN 32 => bit_in_tb <= '0';
                WHEN 33 => bit_in_tb <= '0';
                WHEN 34 => bit_in_tb <= '0';
                WHEN 35 => bit_in_tb <= '1';
                WHEN 36 => bit_in_tb <= '0';
                WHEN 37 => bit_in_tb <= '0';
                WHEN 38 => bit_in_tb <= '1';
                WHEN 39 => bit_in_tb <= '1';
                WHEN 40 => bit_in_tb <= '0';
                WHEN 41 => bit_in_tb <= '1';
                WHEN 42 => bit_in_tb <= '0';
                WHEN 43 => bit_in_tb <= '0';
                WHEN 44 => bit_in_tb <= '0';
                WHEN 45 => bit_in_tb <= '1';
                WHEN 46 => bit_in_tb <= '1';
                WHEN 47 => bit_in_tb <= '0';
                WHEN 48 => bit_in_tb <= '0';
                WHEN 49 => bit_in_tb <= '1';
                WHEN 50 => bit_in_tb <= '0';
                WHEN 51 => bit_in_tb <= '1';
                WHEN 52 => bit_in_tb <= '0';
                WHEN 53 => bit_in_tb <= '1';
                WHEN 54 => bit_in_tb <= '1';
                WHEN 55 => bit_in_tb <= '1';
                WHEN 56 => bit_in_tb <= '1';
                WHEN 57 => bit_in_tb <= '1';
                WHEN 58 => bit_in_tb <= '1';
                WHEN 59 => bit_in_tb <= '1';
                WHEN 60 => bit_in_tb <= '0';
                WHEN 61 => bit_in_tb <= '1';
                WHEN 62 => bit_in_tb <= '1';
                WHEN 63 => bit_in_tb <= '0';
                WHEN 64 => bit_in_tb <= '0';
                WHEN 65 => bit_in_tb <= '1';
                WHEN 66 => bit_in_tb <= '1';
                WHEN 67 => bit_in_tb <= '0';
                WHEN 68 => bit_in_tb <= '0';
                WHEN 69 => bit_in_tb <= '1';
                WHEN 70 => bit_in_tb <= '0';
                WHEN 71 => bit_in_tb <= '0';
                WHEN 72 => bit_in_tb <= '1';
                WHEN 73 => bit_in_tb <= '0';
                WHEN 74 => bit_in_tb <= '0';
                WHEN 75 => bit_in_tb <= '0';
                WHEN 76 => bit_in_tb <= '1';
                WHEN 77 => bit_in_tb <= '1';
                WHEN 78 => bit_in_tb <= '1';
                WHEN 79 => bit_in_tb <= '0';
                WHEN 80 => bit_in_tb <= '1';
                WHEN 81 => bit_in_tb <= '1';
                WHEN 82 => bit_in_tb <= '1';
                WHEN 83 => bit_in_tb <= '0';
                WHEN 84 => bit_in_tb <= '0';
                WHEN 85 => bit_in_tb <= '0';
                WHEN 86 => bit_in_tb <= '1';
                WHEN 87 => bit_in_tb <= '0';
                WHEN 88 => bit_in_tb <= '0';
                WHEN 89 => bit_in_tb <= '0';
                WHEN 90 => bit_in_tb <= '1';
                WHEN 91 => bit_in_tb <= '0';
                WHEN 92 => bit_in_tb <= '0';
                WHEN 93 => bit_in_tb <= '0';
                WHEN 94 => bit_in_tb <= '1';
                WHEN 95 => bit_in_tb <= '1';
                WHEN 96 => bit_in_tb <= '0';
                WHEN 97 => bit_in_tb <= '0';
                WHEN 98 => bit_in_tb <= '1';
                WHEN 99 => bit_in_tb <= '1';
                WHEN 100 => bit_in_tb <= '0';
                WHEN 101 => bit_in_tb <= '1';
                WHEN 102 => bit_in_tb <= '1';
                WHEN 103 => bit_in_tb <= '0';
                WHEN 104 => bit_in_tb <= '0';
                WHEN 105 => bit_in_tb <= '0';
                WHEN 106 => bit_in_tb <= '1';
                WHEN 107 => bit_in_tb <= '0';
                WHEN 108 => bit_in_tb <= '1';
                WHEN 109 => bit_in_tb <= '0';
                WHEN 110 => bit_in_tb <= '0';
                WHEN 111 => bit_in_tb <= '1';
                WHEN 112 => bit_in_tb <= '0';
                WHEN 113 => bit_in_tb <= '0';
                WHEN 114 => bit_in_tb <= '1';
                WHEN 115 => bit_in_tb <= '0';
                WHEN 116 => bit_in_tb <= '0';
                WHEN 117 => bit_in_tb <= '1';
                WHEN 118 => bit_in_tb <= '1';
                WHEN 119 => bit_in_tb <= '1';
                WHEN 120 => bit_in_tb <= '1';
                WHEN 121 => bit_in_tb <= '1';
                WHEN 122 => bit_in_tb <= '0';
                WHEN 123 => bit_in_tb <= '1';
                WHEN 124 => bit_in_tb <= '0';
                WHEN 125 => bit_in_tb <= '0';
                WHEN 126 => bit_in_tb <= '1';
                WHEN 127 => bit_in_tb <= '0';
                WHEN 128 => bit_in_tb <= '1';
                WHEN 129 => bit_in_tb <= '0';
                WHEN 130 => bit_in_tb <= '0';
                WHEN 131 => bit_in_tb <= '1';
                WHEN 132 => bit_in_tb <= '1';
                WHEN 133 => bit_in_tb <= '1';
                WHEN 134 => bit_in_tb <= '0';
                WHEN 135 => bit_in_tb <= '0';
                WHEN 136 => bit_in_tb <= '0';
                WHEN 137 => bit_in_tb <= '0';
                WHEN 138 => bit_in_tb <= '0';
                WHEN 139 => bit_in_tb <= '0';
                WHEN 140 => bit_in_tb <= '0';
                WHEN 141 => bit_in_tb <= '1';
                WHEN 142 => bit_in_tb <= '0';
                WHEN 143 => bit_in_tb <= '1';
                WHEN 144 => bit_in_tb <= '1';
                WHEN 145 => bit_in_tb <= '0';
                WHEN 146 => bit_in_tb <= '1';
                WHEN 147 => bit_in_tb <= '1';
                WHEN 148 => bit_in_tb <= '1';
                WHEN 149 => bit_in_tb <= '1';
                WHEN 150 => bit_in_tb <= '0';
                WHEN 151 => bit_in_tb <= '1';
                WHEN 152 => bit_in_tb <= '0';
                WHEN 153 => bit_in_tb <= '0';
                WHEN 154 => bit_in_tb <= '0';
                WHEN 155 => bit_in_tb <= '0';
                WHEN 156 => bit_in_tb <= '1';
                WHEN 157 => bit_in_tb <= '0';
                WHEN 158 => bit_in_tb <= '0';
                WHEN 159 => bit_in_tb <= '0';
                WHEN 160 => bit_in_tb <= '1';
                WHEN 161 => bit_in_tb <= '1';
                WHEN 162 => bit_in_tb <= '0';
                WHEN 163 => bit_in_tb <= '0';
                WHEN 164 => bit_in_tb <= '0';
                WHEN 165 => bit_in_tb <= '0';
                WHEN 166 => bit_in_tb <= '0';
                WHEN 167 => bit_in_tb <= '0';
                WHEN 168 => bit_in_tb <= '1';
                WHEN 169 => bit_in_tb <= '0';
                WHEN 170 => bit_in_tb <= '0';
                WHEN 171 => bit_in_tb <= '0';
                WHEN 172 => bit_in_tb <= '1';
                WHEN 173 => bit_in_tb <= '1';
                WHEN 174 => bit_in_tb <= '1';
                WHEN 175 => bit_in_tb <= '1';
                WHEN 176 => bit_in_tb <= '1';
                WHEN 177 => bit_in_tb <= '1';
                WHEN 178 => bit_in_tb <= '1';
                WHEN 179 => bit_in_tb <= '1';
                WHEN 180 => bit_in_tb <= '1';
                WHEN 181 => bit_in_tb <= '1';
                WHEN 182 => bit_in_tb <= '0';
                WHEN 183 => bit_in_tb <= '1';
                WHEN 184 => bit_in_tb <= '0';
                WHEN 185 => bit_in_tb <= '0';
                WHEN 186 => bit_in_tb <= '0';
                WHEN 187 => bit_in_tb <= '0';
                WHEN 188 => bit_in_tb <= '1';
                WHEN 189 => bit_in_tb <= '1';
                WHEN 190 => bit_in_tb <= '1';
                WHEN 191 => bit_in_tb <= '0';
                WHEN 192 => bit_in_tb <= '1';
                WHEN 193 => bit_in_tb <= '0';
                WHEN 194 => bit_in_tb <= '1';
                WHEN 195 => bit_in_tb <= '1';
                WHEN 196 => bit_in_tb <= '1';
                WHEN 197 => bit_in_tb <= '0';
                WHEN 198 => bit_in_tb <= '0';
                WHEN 199 => bit_in_tb <= '0';
                WHEN 200 => bit_in_tb <= '0';
                WHEN 201 => bit_in_tb <= '0';
                WHEN 202 => bit_in_tb <= '0';
                WHEN 203 => bit_in_tb <= '1';
                WHEN 204 => bit_in_tb <= '1';
                WHEN 205 => bit_in_tb <= '0';
                WHEN 206 => bit_in_tb <= '1';
                WHEN 207 => bit_in_tb <= '1';
                WHEN 208 => bit_in_tb <= '0';
                WHEN 209 => bit_in_tb <= '0';
                WHEN 210 => bit_in_tb <= '1';
                WHEN 211 => bit_in_tb <= '1';
                WHEN 212 => bit_in_tb <= '1';
                WHEN 213 => bit_in_tb <= '0';
                WHEN 214 => bit_in_tb <= '0';
                WHEN 215 => bit_in_tb <= '1';
                WHEN 216 => bit_in_tb <= '0';
                WHEN 217 => bit_in_tb <= '0';
                WHEN 218 => bit_in_tb <= '1';
                WHEN 219 => bit_in_tb <= '1';
                WHEN 220 => bit_in_tb <= '0';
                WHEN 221 => bit_in_tb <= '1';
                WHEN 222 => bit_in_tb <= '0';
                WHEN 223 => bit_in_tb <= '1';
                WHEN 224 => bit_in_tb <= '1';
                WHEN 225 => bit_in_tb <= '1';
                WHEN 226 => bit_in_tb <= '0';
                WHEN 227 => bit_in_tb <= '0';
                WHEN 228 => bit_in_tb <= '0';
                WHEN 229 => bit_in_tb <= '1';
                WHEN 230 => bit_in_tb <= '1';
                WHEN 231 => bit_in_tb <= '0';
                WHEN 232 => bit_in_tb <= '0';
                WHEN 233 => bit_in_tb <= '0';
                WHEN 234 => bit_in_tb <= '1';
                WHEN 235 => bit_in_tb <= '1';
                WHEN 236 => bit_in_tb <= '0';
                WHEN 237 => bit_in_tb <= '0';
                WHEN 238 => bit_in_tb <= '0';
                WHEN 239 => bit_in_tb <= '1';
                WHEN 240 => bit_in_tb <= '1';
                WHEN 241 => bit_in_tb <= '1';
                WHEN 242 => bit_in_tb <= '0';
                WHEN 243 => bit_in_tb <= '1';
                WHEN 244 => bit_in_tb <= '0';
                WHEN 245 => bit_in_tb <= '1';
                WHEN 246 => bit_in_tb <= '0';
                WHEN 247 => bit_in_tb <= '0';
                WHEN 248 => bit_in_tb <= '0';
                WHEN 249 => bit_in_tb <= '1';
                WHEN 250 => bit_in_tb <= '0';
                WHEN 251 => bit_in_tb <= '0';
                WHEN 252 => bit_in_tb <= '0';
                WHEN 253 => bit_in_tb <= '1';
                WHEN 254 => bit_in_tb <= '0';
                WHEN 255 => bit_in_tb <= '0';
                WHEN 256 => bit_in_tb <= '0';
                WHEN 257 => bit_in_tb <= '0';
                WHEN 258 => bit_in_tb <= '0';
                WHEN 259 => bit_in_tb <= '1';
                WHEN 260 => bit_in_tb <= '0';
                WHEN 261 => bit_in_tb <= '0';
                WHEN 262 => bit_in_tb <= '1';
                WHEN 263 => bit_in_tb <= '0';
                WHEN 264 => bit_in_tb <= '0';
                WHEN 265 => bit_in_tb <= '1';
                WHEN 266 => bit_in_tb <= '1';
                WHEN 267 => bit_in_tb <= '0';
                WHEN 268 => bit_in_tb <= '0';
                WHEN 269 => bit_in_tb <= '0';
                WHEN 270 => bit_in_tb <= '0';
                WHEN 271 => bit_in_tb <= '1';
                WHEN 272 => bit_in_tb <= '0';
                WHEN 273 => bit_in_tb <= '0';
                WHEN 274 => bit_in_tb <= '0';
                WHEN 275 => bit_in_tb <= '1';
                WHEN 276 => bit_in_tb <= '1';
                WHEN 277 => bit_in_tb <= '0';
                WHEN 278 => bit_in_tb <= '1';
                WHEN 279 => bit_in_tb <= '1';
                WHEN 280 => bit_in_tb <= '0';
                WHEN 281 => bit_in_tb <= '1';
                WHEN 282 => bit_in_tb <= '0';
                WHEN 283 => bit_in_tb <= '1';
                WHEN 284 => bit_in_tb <= '1';
                WHEN 285 => bit_in_tb <= '1';
                WHEN 286 => bit_in_tb <= '1';
                WHEN 287 => bit_in_tb <= '1';
                WHEN 288 => bit_in_tb <= '0';
                WHEN 289 => bit_in_tb <= '0';
                WHEN 290 => bit_in_tb <= '1';
                WHEN 291 => bit_in_tb <= '1';
                WHEN 292 => bit_in_tb <= '0';
                WHEN 293 => bit_in_tb <= '1';
                WHEN 294 => bit_in_tb <= '1';
                WHEN 295 => bit_in_tb <= '0';
                WHEN 296 => bit_in_tb <= '0';
                WHEN 297 => bit_in_tb <= '1';
                WHEN 298 => bit_in_tb <= '0';
                WHEN 299 => bit_in_tb <= '1';
                WHEN 300 => bit_in_tb <= '0';
                WHEN 301 => bit_in_tb <= '0';
                WHEN 302 => bit_in_tb <= '0';
                WHEN 303 => bit_in_tb <= '1';
                WHEN 304 => bit_in_tb <= '0';
                WHEN 305 => bit_in_tb <= '0';
                WHEN 306 => bit_in_tb <= '1';
                WHEN 307 => bit_in_tb <= '1';
                WHEN 308 => bit_in_tb <= '0';
                WHEN 309 => bit_in_tb <= '1';
                WHEN 310 => bit_in_tb <= '1';
                WHEN 311 => bit_in_tb <= '1';
                WHEN 312 => bit_in_tb <= '0';
                WHEN 313 => bit_in_tb <= '0';
                WHEN 314 => bit_in_tb <= '0';
                WHEN 315 => bit_in_tb <= '1';
                WHEN 316 => bit_in_tb <= '1';
                WHEN 317 => bit_in_tb <= '1';
                WHEN 318 => bit_in_tb <= '0';
                WHEN 319 => bit_in_tb <= '0';
                WHEN 320 => bit_in_tb <= '0';
                WHEN 321 => bit_in_tb <= '1';
                WHEN 322 => bit_in_tb <= '1';
                WHEN 323 => bit_in_tb <= '0';
                WHEN 324 => bit_in_tb <= '0';
                WHEN 325 => bit_in_tb <= '1';
                WHEN 326 => bit_in_tb <= '1';
                WHEN 327 => bit_in_tb <= '0';
                WHEN 328 => bit_in_tb <= '0';
                WHEN 329 => bit_in_tb <= '0';
                WHEN 330 => bit_in_tb <= '1';
                WHEN 331 => bit_in_tb <= '0';
                WHEN 332 => bit_in_tb <= '0';
                WHEN 333 => bit_in_tb <= '0';
                WHEN 334 => bit_in_tb <= '1';
                WHEN 335 => bit_in_tb <= '1';
                WHEN 336 => bit_in_tb <= '1';
                WHEN 337 => bit_in_tb <= '1';
                WHEN 338 => bit_in_tb <= '1';
                WHEN 339 => bit_in_tb <= '0';
                WHEN 340 => bit_in_tb <= '0';
                WHEN 341 => bit_in_tb <= '0';
                WHEN 342 => bit_in_tb <= '1';
                WHEN 343 => bit_in_tb <= '0';
                WHEN 344 => bit_in_tb <= '1';
                WHEN 345 => bit_in_tb <= '1';
                WHEN 346 => bit_in_tb <= '1';
                WHEN 347 => bit_in_tb <= '1';
                WHEN 348 => bit_in_tb <= '1';
                WHEN 349 => bit_in_tb <= '0';
                WHEN 350 => bit_in_tb <= '1';
                WHEN 351 => bit_in_tb <= '0';
                WHEN 352 => bit_in_tb <= '1';
                WHEN 353 => bit_in_tb <= '0';
                WHEN 354 => bit_in_tb <= '0';
                WHEN 355 => bit_in_tb <= '1';
                WHEN 356 => bit_in_tb <= '0';
                WHEN 357 => bit_in_tb <= '1';
                WHEN 358 => bit_in_tb <= '1';
                WHEN 359 => bit_in_tb <= '0';
                WHEN 360 => bit_in_tb <= '1';
                WHEN 361 => bit_in_tb <= '0';
                WHEN 362 => bit_in_tb <= '0';
                WHEN 363 => bit_in_tb <= '1';
                WHEN 364 => bit_in_tb <= '1';
                WHEN 365 => bit_in_tb <= '1';
                WHEN 366 => bit_in_tb <= '0';
                WHEN 367 => bit_in_tb <= '1';
                WHEN 368 => bit_in_tb <= '0';
                WHEN 369 => bit_in_tb <= '0';
                WHEN 370 => bit_in_tb <= '1';
                WHEN 371 => bit_in_tb <= '0';
                WHEN 372 => bit_in_tb <= '0';
                WHEN 373 => bit_in_tb <= '0';
                WHEN 374 => bit_in_tb <= '0';
                WHEN 375 => bit_in_tb <= '0';
                WHEN 376 => bit_in_tb <= '1';
                WHEN 377 => bit_in_tb <= '0';
                WHEN 378 => bit_in_tb <= '1';
                WHEN 379 => bit_in_tb <= '0';
                WHEN 380 => bit_in_tb <= '1';
                WHEN 381 => bit_in_tb <= '0';
                WHEN 382 => bit_in_tb <= '0';
                WHEN 383 => bit_in_tb <= '0';
                WHEN 384 => bit_in_tb <= '1';
                WHEN 385 => bit_in_tb <= '0';
                WHEN 386 => bit_in_tb <= '1';
                WHEN 387 => bit_in_tb <= '1';
                WHEN 388 => bit_in_tb <= '1';
                WHEN 389 => bit_in_tb <= '1';
                WHEN 390 => bit_in_tb <= '1';
                WHEN 391 => bit_in_tb <= '1';
                WHEN 392 => bit_in_tb <= '1';
                WHEN 393 => bit_in_tb <= '0';
                WHEN 394 => bit_in_tb <= '1';
                WHEN 395 => bit_in_tb <= '1';
                WHEN 396 => bit_in_tb <= '0';
                WHEN 397 => bit_in_tb <= '1';
                WHEN 398 => bit_in_tb <= '0';
                WHEN 399 => bit_in_tb <= '1';
                WHEN 400 => bit_in_tb <= '0';
                WHEN 401 => bit_in_tb <= '0';
                WHEN 402 => bit_in_tb <= '0';
                WHEN 403 => bit_in_tb <= '0';
                WHEN 404 => bit_in_tb <= '1';
                WHEN 405 => bit_in_tb <= '0';
                WHEN 406 => bit_in_tb <= '0';
                WHEN 407 => bit_in_tb <= '1';
                WHEN 408 => bit_in_tb <= '1';
                WHEN 409 => bit_in_tb <= '1';
                WHEN 410 => bit_in_tb <= '1';
                WHEN 411 => bit_in_tb <= '1';
                WHEN 412 => bit_in_tb <= '1';
                WHEN 413 => bit_in_tb <= '0';
                WHEN 414 => bit_in_tb <= '1';
                WHEN 415 => bit_in_tb <= '0';
                WHEN 416 => bit_in_tb <= '1';
                WHEN 417 => bit_in_tb <= '0';
                WHEN 418 => bit_in_tb <= '1';
                WHEN 419 => bit_in_tb <= '0';
                WHEN 420 => bit_in_tb <= '0';
                WHEN 421 => bit_in_tb <= '0';
                WHEN 422 => bit_in_tb <= '1';
                WHEN 423 => bit_in_tb <= '1';
                WHEN 424 => bit_in_tb <= '1';
                WHEN 425 => bit_in_tb <= '0';
                WHEN 426 => bit_in_tb <= '1';
                WHEN 427 => bit_in_tb <= '0';
                WHEN 428 => bit_in_tb <= '0';
                WHEN 429 => bit_in_tb <= '1';
                WHEN 430 => bit_in_tb <= '0';
                WHEN 431 => bit_in_tb <= '0';
                WHEN 432 => bit_in_tb <= '0';
                WHEN 433 => bit_in_tb <= '0';
                WHEN 434 => bit_in_tb <= '0';
                WHEN 435 => bit_in_tb <= '1';
                WHEN 436 => bit_in_tb <= '0';
                WHEN 437 => bit_in_tb <= '1';
                WHEN 438 => bit_in_tb <= '0';
                WHEN 439 => bit_in_tb <= '0';
                WHEN 440 => bit_in_tb <= '1';
                WHEN 441 => bit_in_tb <= '1';
                WHEN 442 => bit_in_tb <= '1';
                WHEN 443 => bit_in_tb <= '1';
                WHEN 444 => bit_in_tb <= '1';
                WHEN 445 => bit_in_tb <= '1';
                WHEN 446 => bit_in_tb <= '1';
                WHEN 447 => bit_in_tb <= '1';
                WHEN 448 => bit_in_tb <= '0';
                WHEN 449 => bit_in_tb <= '1';
                WHEN 450 => bit_in_tb <= '1';
                WHEN 451 => bit_in_tb <= '1';
                WHEN 452 => bit_in_tb <= '1';
                WHEN 453 => bit_in_tb <= '1';
                WHEN 454 => bit_in_tb <= '1';
                WHEN 455 => bit_in_tb <= '0';
                WHEN 456 => bit_in_tb <= '0';
                WHEN 457 => bit_in_tb <= '1';
                WHEN 458 => bit_in_tb <= '0';
                WHEN 459 => bit_in_tb <= '1';
                WHEN 460 => bit_in_tb <= '0';
                WHEN 461 => bit_in_tb <= '1';
                WHEN 462 => bit_in_tb <= '1';
                WHEN 463 => bit_in_tb <= '1';
                WHEN 464 => bit_in_tb <= '1';
                WHEN 465 => bit_in_tb <= '1';
                WHEN 466 => bit_in_tb <= '0';
                WHEN 467 => bit_in_tb <= '0';
                WHEN 468 => bit_in_tb <= '0';
                WHEN 469 => bit_in_tb <= '1';
                WHEN 470 => bit_in_tb <= '0';
                WHEN 471 => bit_in_tb <= '1';
                WHEN 472 => bit_in_tb <= '1';
                WHEN 473 => bit_in_tb <= '1';
                WHEN 474 => bit_in_tb <= '0';
                WHEN 475 => bit_in_tb <= '0';
                WHEN 476 => bit_in_tb <= '1';
                WHEN 477 => bit_in_tb <= '1';
                WHEN 478 => bit_in_tb <= '0';
                WHEN 479 => bit_in_tb <= '0';
                WHEN 480 => bit_in_tb <= '1';
                WHEN 481 => bit_in_tb <= '1';
                WHEN 482 => bit_in_tb <= '0';
                WHEN 483 => bit_in_tb <= '1';
                WHEN 484 => bit_in_tb <= '1';
                WHEN 485 => bit_in_tb <= '1';
                WHEN 486 => bit_in_tb <= '1';
                WHEN 487 => bit_in_tb <= '1';
                WHEN 488 => bit_in_tb <= '0';
                WHEN 489 => bit_in_tb <= '0';
                WHEN 490 => bit_in_tb <= '0';
                WHEN 491 => bit_in_tb <= '1';
                WHEN 492 => bit_in_tb <= '0';
                WHEN 493 => bit_in_tb <= '0';
                WHEN 494 => bit_in_tb <= '0';
                WHEN 495 => bit_in_tb <= '0';
                WHEN 496 => bit_in_tb <= '0';
                WHEN 497 => bit_in_tb <= '1';
                WHEN 498 => bit_in_tb <= '0';
                WHEN 499 => bit_in_tb <= '0';
                WHEN 500 => bit_in_tb <= '0';
                WHEN 501 => bit_in_tb <= '0';
                WHEN 502 => bit_in_tb <= '1';
                WHEN 503 => bit_in_tb <= '0';
                WHEN 504 => bit_in_tb <= '0';
                WHEN 505 => bit_in_tb <= '0';
                WHEN 506 => bit_in_tb <= '0';
                WHEN 507 => bit_in_tb <= '1';
                WHEN 508 => bit_in_tb <= '0';
                WHEN 509 => bit_in_tb <= '0';
                WHEN 510 => bit_in_tb <= '1';
                WHEN 511 => bit_in_tb <= '1';
                WHEN 512 => bit_in_tb <= '0';
                WHEN 513 => bit_in_tb <= '1';
                WHEN 514 => bit_in_tb <= '1';
                WHEN 515 => bit_in_tb <= '0';
                WHEN 516 => bit_in_tb <= '0';
                WHEN 517 => bit_in_tb <= '0';
                WHEN 518 => bit_in_tb <= '0';
                WHEN 519 => bit_in_tb <= '0';
                WHEN 520 => bit_in_tb <= '1';
                WHEN 521 => bit_in_tb <= '1';
                WHEN 522 => bit_in_tb <= '1';
                WHEN 523 => bit_in_tb <= '1';
                WHEN 524 => bit_in_tb <= '1';
                WHEN 525 => bit_in_tb <= '1';
                WHEN 526 => bit_in_tb <= '1';
                WHEN 527 => bit_in_tb <= '1';
                WHEN 528 => bit_in_tb <= '0';
                WHEN 529 => bit_in_tb <= '0';
                WHEN 530 => bit_in_tb <= '0';
                WHEN 531 => bit_in_tb <= '1';
                WHEN 532 => bit_in_tb <= '0';
                WHEN 533 => bit_in_tb <= '1';
                WHEN 534 => bit_in_tb <= '1';
                WHEN 535 => bit_in_tb <= '1';
                WHEN 536 => bit_in_tb <= '1';
                WHEN 537 => bit_in_tb <= '0';
                WHEN 538 => bit_in_tb <= '1';
                WHEN 539 => bit_in_tb <= '1';
                WHEN 540 => bit_in_tb <= '1';
                WHEN 541 => bit_in_tb <= '0';
                WHEN 542 => bit_in_tb <= '0';
                WHEN 543 => bit_in_tb <= '1';
                WHEN 544 => bit_in_tb <= '1';
                WHEN 545 => bit_in_tb <= '0';
                WHEN 546 => bit_in_tb <= '0';
                WHEN 547 => bit_in_tb <= '0';
                WHEN 548 => bit_in_tb <= '1';
                WHEN 549 => bit_in_tb <= '1';
                WHEN 550 => bit_in_tb <= '1';
                WHEN 551 => bit_in_tb <= '0';
                WHEN 552 => bit_in_tb <= '1';
                WHEN 553 => bit_in_tb <= '1';
                WHEN 554 => bit_in_tb <= '1';
                WHEN 555 => bit_in_tb <= '1';
                WHEN 556 => bit_in_tb <= '1';
                WHEN 557 => bit_in_tb <= '1';
                WHEN 558 => bit_in_tb <= '1';
                WHEN 559 => bit_in_tb <= '0';
                WHEN 560 => bit_in_tb <= '1';
                WHEN 561 => bit_in_tb <= '1';
                WHEN 562 => bit_in_tb <= '1';
                WHEN 563 => bit_in_tb <= '1';
                WHEN 564 => bit_in_tb <= '0';
                WHEN 565 => bit_in_tb <= '0';
                WHEN 566 => bit_in_tb <= '0';
                WHEN 567 => bit_in_tb <= '0';
                WHEN 568 => bit_in_tb <= '1';
                WHEN 569 => bit_in_tb <= '1';
                WHEN 570 => bit_in_tb <= '0';
                WHEN 571 => bit_in_tb <= '0';
                WHEN 572 => bit_in_tb <= '0';
                WHEN 573 => bit_in_tb <= '1';
                WHEN 574 => bit_in_tb <= '0';
                WHEN 575 => bit_in_tb <= '1';
                WHEN 576 => bit_in_tb <= '0';
                WHEN 577 => bit_in_tb <= '0';
                WHEN 578 => bit_in_tb <= '1';
                WHEN 579 => bit_in_tb <= '0';
                WHEN 580 => bit_in_tb <= '1';
                WHEN 581 => bit_in_tb <= '0';
                WHEN 582 => bit_in_tb <= '1';
                WHEN 583 => bit_in_tb <= '1';
                WHEN 584 => bit_in_tb <= '0';
                WHEN 585 => bit_in_tb <= '0';
                WHEN 586 => bit_in_tb <= '1';
                WHEN 587 => bit_in_tb <= '0';
                WHEN 588 => bit_in_tb <= '0';
                WHEN 589 => bit_in_tb <= '1';
                WHEN 590 => bit_in_tb <= '0';
                WHEN 591 => bit_in_tb <= '0';
                WHEN 592 => bit_in_tb <= '0';
                WHEN 593 => bit_in_tb <= '1';
                WHEN 594 => bit_in_tb <= '1';
                WHEN 595 => bit_in_tb <= '0';
                WHEN 596 => bit_in_tb <= '1';
                WHEN 597 => bit_in_tb <= '0';
                WHEN 598 => bit_in_tb <= '1';
                WHEN 599 => bit_in_tb <= '0';
                WHEN 600 => bit_in_tb <= '0';
                WHEN 601 => bit_in_tb <= '0';
                WHEN 602 => bit_in_tb <= '1';
                WHEN 603 => bit_in_tb <= '0';
                WHEN 604 => bit_in_tb <= '1';
                WHEN 605 => bit_in_tb <= '0';
                WHEN 606 => bit_in_tb <= '1';
                WHEN 607 => bit_in_tb <= '1';
                WHEN 608 => bit_in_tb <= '0';
                WHEN 609 => bit_in_tb <= '0';
                WHEN 610 => bit_in_tb <= '1';
                WHEN 611 => bit_in_tb <= '0';
                WHEN 612 => bit_in_tb <= '1';
                WHEN 613 => bit_in_tb <= '1';
                WHEN 614 => bit_in_tb <= '0';
                WHEN 615 => bit_in_tb <= '1';
                WHEN 616 => bit_in_tb <= '1';
                WHEN 617 => bit_in_tb <= '1';
                WHEN 618 => bit_in_tb <= '1';
                WHEN 619 => bit_in_tb <= '0';
                WHEN 620 => bit_in_tb <= '1';
                WHEN 621 => bit_in_tb <= '0';
                WHEN 622 => bit_in_tb <= '0';
                WHEN 623 => bit_in_tb <= '1';
                WHEN 624 => bit_in_tb <= '1';
                WHEN 625 => bit_in_tb <= '0';
                WHEN 626 => bit_in_tb <= '0';
                WHEN 627 => bit_in_tb <= '0';
                WHEN 628 => bit_in_tb <= '1';
                WHEN 629 => bit_in_tb <= '1';
                WHEN 630 => bit_in_tb <= '0';
                WHEN 631 => bit_in_tb <= '1';
                WHEN 632 => bit_in_tb <= '1';
                WHEN 633 => bit_in_tb <= '0';
                WHEN 634 => bit_in_tb <= '1';
                WHEN 635 => bit_in_tb <= '1';
                WHEN 636 => bit_in_tb <= '1';
                WHEN 637 => bit_in_tb <= '1';
                WHEN 638 => bit_in_tb <= '1';
                WHEN 639 => bit_in_tb <= '0';
                WHEN 640 => bit_in_tb <= '0';
                WHEN 641 => bit_in_tb <= '1';
                WHEN 642 => bit_in_tb <= '0';
                WHEN 643 => bit_in_tb <= '1';
                WHEN 644 => bit_in_tb <= '0';
                WHEN 645 => bit_in_tb <= '1';
                WHEN 646 => bit_in_tb <= '0';
                WHEN 647 => bit_in_tb <= '0';
                WHEN 648 => bit_in_tb <= '0';
                WHEN 649 => bit_in_tb <= '0';
                WHEN 650 => bit_in_tb <= '0';
                WHEN 651 => bit_in_tb <= '1';
                WHEN 652 => bit_in_tb <= '1';
                WHEN 653 => bit_in_tb <= '1';
                WHEN 654 => bit_in_tb <= '0';
                WHEN 655 => bit_in_tb <= '0';
                WHEN 656 => bit_in_tb <= '1';
                WHEN 657 => bit_in_tb <= '0';
                WHEN 658 => bit_in_tb <= '0';
                WHEN 659 => bit_in_tb <= '0';
                WHEN 660 => bit_in_tb <= '1';
                WHEN 661 => bit_in_tb <= '1';
                WHEN 662 => bit_in_tb <= '0';
                WHEN 663 => bit_in_tb <= '1';
                WHEN 664 => bit_in_tb <= '1';
                WHEN 665 => bit_in_tb <= '1';
                WHEN 666 => bit_in_tb <= '0';
                WHEN 667 => bit_in_tb <= '0';
                WHEN 668 => bit_in_tb <= '0';
                WHEN 669 => bit_in_tb <= '1';
                WHEN 670 => bit_in_tb <= '1';
                WHEN 671 => bit_in_tb <= '1';
                WHEN 672 => bit_in_tb <= '0';
                WHEN 673 => bit_in_tb <= '1';
                WHEN 674 => bit_in_tb <= '1';
                WHEN 675 => bit_in_tb <= '0';
                WHEN 676 => bit_in_tb <= '1';
                WHEN 677 => bit_in_tb <= '1';
                WHEN 678 => bit_in_tb <= '1';
                WHEN 679 => bit_in_tb <= '0';
                WHEN 680 => bit_in_tb <= '0';
                WHEN 681 => bit_in_tb <= '1';
                WHEN 682 => bit_in_tb <= '1';
                WHEN 683 => bit_in_tb <= '0';
                WHEN 684 => bit_in_tb <= '0';
                WHEN 685 => bit_in_tb <= '0';
                WHEN 686 => bit_in_tb <= '1';
                WHEN 687 => bit_in_tb <= '0';
                WHEN 688 => bit_in_tb <= '0';
                WHEN 689 => bit_in_tb <= '1';
                WHEN 690 => bit_in_tb <= '0';
                WHEN 691 => bit_in_tb <= '1';
                WHEN 692 => bit_in_tb <= '1';
                WHEN 693 => bit_in_tb <= '0';
                WHEN 694 => bit_in_tb <= '0';
                WHEN 695 => bit_in_tb <= '0';
                WHEN 696 => bit_in_tb <= '0';
                WHEN 697 => bit_in_tb <= '1';
                WHEN 698 => bit_in_tb <= '1';
                WHEN 699 => bit_in_tb <= '1';
                WHEN 700 => bit_in_tb <= '0';
                WHEN 701 => bit_in_tb <= '1';
                WHEN 702 => bit_in_tb <= '1';
                WHEN 703 => bit_in_tb <= '0';
                WHEN 704 => bit_in_tb <= '1';
                WHEN 705 => bit_in_tb <= '0';
                WHEN 706 => bit_in_tb <= '0';
                WHEN 707 => bit_in_tb <= '0';
                WHEN 708 => bit_in_tb <= '0';
                WHEN 709 => bit_in_tb <= '0';
                WHEN 710 => bit_in_tb <= '0';
                WHEN 711 => bit_in_tb <= '0';
                WHEN 712 => bit_in_tb <= '0';
                WHEN 713 => bit_in_tb <= '1';
                WHEN 714 => bit_in_tb <= '1';
                WHEN 715 => bit_in_tb <= '1';
                WHEN 716 => bit_in_tb <= '0';
                WHEN 717 => bit_in_tb <= '0';
                WHEN 718 => bit_in_tb <= '1';
                WHEN 719 => bit_in_tb <= '1';
                WHEN 720 => bit_in_tb <= '1';
                WHEN 721 => bit_in_tb <= '0';
                WHEN 722 => bit_in_tb <= '0';
                WHEN 723 => bit_in_tb <= '0';
                WHEN 724 => bit_in_tb <= '0';
                WHEN 725 => bit_in_tb <= '0';
                WHEN 726 => bit_in_tb <= '1';
                WHEN 727 => bit_in_tb <= '1';
                WHEN 728 => bit_in_tb <= '1';
                WHEN 729 => bit_in_tb <= '0';
                WHEN 730 => bit_in_tb <= '1';
                WHEN 731 => bit_in_tb <= '0';
                WHEN 732 => bit_in_tb <= '0';
                WHEN 733 => bit_in_tb <= '1';
                WHEN 734 => bit_in_tb <= '0';
                WHEN 735 => bit_in_tb <= '0';
                WHEN 736 => bit_in_tb <= '0';
                WHEN 737 => bit_in_tb <= '0';
                WHEN 738 => bit_in_tb <= '1';
                WHEN 739 => bit_in_tb <= '1';
                WHEN 740 => bit_in_tb <= '0';
                WHEN 741 => bit_in_tb <= '1';
                WHEN 742 => bit_in_tb <= '1';
                WHEN 743 => bit_in_tb <= '0';
                WHEN 744 => bit_in_tb <= '0';
                WHEN 745 => bit_in_tb <= '1';
                WHEN 746 => bit_in_tb <= '1';
                WHEN 747 => bit_in_tb <= '0';
                WHEN 748 => bit_in_tb <= '0';
                WHEN 749 => bit_in_tb <= '1';
                WHEN 750 => bit_in_tb <= '0';
                WHEN 751 => bit_in_tb <= '1';
                WHEN 752 => bit_in_tb <= '1';
                WHEN 753 => bit_in_tb <= '0';
                WHEN 754 => bit_in_tb <= '1';
                WHEN 755 => bit_in_tb <= '0';
                WHEN 756 => bit_in_tb <= '0';
                WHEN 757 => bit_in_tb <= '0';
                WHEN 758 => bit_in_tb <= '0';
                WHEN 759 => bit_in_tb <= '1';
                WHEN 760 => bit_in_tb <= '0';
                WHEN 761 => bit_in_tb <= '0';
                WHEN 762 => bit_in_tb <= '1';
                WHEN 763 => bit_in_tb <= '1';
                WHEN 764 => bit_in_tb <= '0';
                WHEN 765 => bit_in_tb <= '1';
                WHEN 766 => bit_in_tb <= '1';
                WHEN 767 => bit_in_tb <= '0';
                WHEN 768 => bit_in_tb <= '1';
                WHEN 769 => bit_in_tb <= '1';
                WHEN 770 => bit_in_tb <= '1';
                WHEN 771 => bit_in_tb <= '1';
                WHEN 772 => bit_in_tb <= '0';
                WHEN 773 => bit_in_tb <= '1';
                WHEN 774 => bit_in_tb <= '1';
                WHEN 775 => bit_in_tb <= '1';
                WHEN 776 => bit_in_tb <= '1';
                WHEN 777 => bit_in_tb <= '1';
                WHEN 778 => bit_in_tb <= '1';
                WHEN 779 => bit_in_tb <= '0';
                WHEN 780 => bit_in_tb <= '0';
                WHEN 781 => bit_in_tb <= '0';
                WHEN 782 => bit_in_tb <= '1';
                WHEN 783 => bit_in_tb <= '0';
                WHEN 784 => bit_in_tb <= '1';
                WHEN 785 => bit_in_tb <= '0';
                WHEN 786 => bit_in_tb <= '0';
                WHEN 787 => bit_in_tb <= '1';
                WHEN 788 => bit_in_tb <= '1';
                WHEN 789 => bit_in_tb <= '0';
                WHEN 790 => bit_in_tb <= '1';
                WHEN 791 => bit_in_tb <= '0';
                WHEN 792 => bit_in_tb <= '0';
                WHEN 793 => bit_in_tb <= '0';
                WHEN 794 => bit_in_tb <= '0';
                WHEN 795 => bit_in_tb <= '1';
                WHEN 796 => bit_in_tb <= '0';
                WHEN 797 => bit_in_tb <= '0';
                WHEN 798 => bit_in_tb <= '0';
                WHEN 799 => bit_in_tb <= '1';
                WHEN 800 => bit_in_tb <= '0';
                WHEN 801 => bit_in_tb <= '0';
                WHEN 802 => bit_in_tb <= '1';
                WHEN 803 => bit_in_tb <= '1';
                WHEN 804 => bit_in_tb <= '1';
                WHEN 805 => bit_in_tb <= '0';
                WHEN 806 => bit_in_tb <= '0';
                WHEN 807 => bit_in_tb <= '0';
                WHEN 808 => bit_in_tb <= '0';
                WHEN 809 => bit_in_tb <= '1';
                WHEN 810 => bit_in_tb <= '0';
                WHEN 811 => bit_in_tb <= '0';
                WHEN 812 => bit_in_tb <= '0';
                WHEN 813 => bit_in_tb <= '1';
                WHEN 814 => bit_in_tb <= '1';
                WHEN 815 => bit_in_tb <= '1';
                WHEN 816 => bit_in_tb <= '0';
                WHEN 817 => bit_in_tb <= '1';
                WHEN 818 => bit_in_tb <= '1';
                WHEN 819 => bit_in_tb <= '0';
                WHEN 820 => bit_in_tb <= '1';
                WHEN 821 => bit_in_tb <= '0';
                WHEN 822 => bit_in_tb <= '1';
                WHEN 823 => bit_in_tb <= '1';
                WHEN 824 => bit_in_tb <= '1';
                WHEN 825 => bit_in_tb <= '1';
                WHEN 826 => bit_in_tb <= '0';
                WHEN 827 => bit_in_tb <= '1';
                WHEN 828 => bit_in_tb <= '1';
                WHEN 829 => bit_in_tb <= '0';
                WHEN 830 => bit_in_tb <= '0';
                WHEN 831 => bit_in_tb <= '1';
                WHEN 832 => bit_in_tb <= '1';
                WHEN 833 => bit_in_tb <= '0';
                WHEN 834 => bit_in_tb <= '0';
                WHEN 835 => bit_in_tb <= '0';
                WHEN 836 => bit_in_tb <= '1';
                WHEN 837 => bit_in_tb <= '1';
                WHEN 838 => bit_in_tb <= '1';
                WHEN 839 => bit_in_tb <= '0';
                WHEN 840 => bit_in_tb <= '1';
                WHEN 841 => bit_in_tb <= '0';
                WHEN 842 => bit_in_tb <= '0';
                WHEN 843 => bit_in_tb <= '1';
                WHEN 844 => bit_in_tb <= '1';
                WHEN 845 => bit_in_tb <= '0';
                WHEN 846 => bit_in_tb <= '0';
                WHEN 847 => bit_in_tb <= '1';
                WHEN 848 => bit_in_tb <= '0';
                WHEN 849 => bit_in_tb <= '0';
                WHEN 850 => bit_in_tb <= '0';
                WHEN 851 => bit_in_tb <= '1';
                WHEN 852 => bit_in_tb <= '0';
                WHEN 853 => bit_in_tb <= '0';
                WHEN 854 => bit_in_tb <= '1';
                WHEN 855 => bit_in_tb <= '1';
                WHEN 856 => bit_in_tb <= '1';
                WHEN 857 => bit_in_tb <= '0';
                WHEN 858 => bit_in_tb <= '1';
                WHEN 859 => bit_in_tb <= '0';
                WHEN 860 => bit_in_tb <= '1';
                WHEN 861 => bit_in_tb <= '0';
                WHEN 862 => bit_in_tb <= '0';
                WHEN 863 => bit_in_tb <= '1';
                WHEN 864 => bit_in_tb <= '1';
                WHEN 865 => bit_in_tb <= '1';
                WHEN 866 => bit_in_tb <= '1';
                WHEN 867 => bit_in_tb <= '0';
                WHEN 868 => bit_in_tb <= '0';
                WHEN 869 => bit_in_tb <= '0';
                WHEN 870 => bit_in_tb <= '0';
                WHEN 871 => bit_in_tb <= '1';
                WHEN 872 => bit_in_tb <= '1';
                WHEN 873 => bit_in_tb <= '0';
                WHEN 874 => bit_in_tb <= '1';
                WHEN 875 => bit_in_tb <= '0';
                WHEN 876 => bit_in_tb <= '0';
                WHEN 877 => bit_in_tb <= '0';
                WHEN 878 => bit_in_tb <= '0';
                WHEN 879 => bit_in_tb <= '1';
                WHEN 880 => bit_in_tb <= '0';
                WHEN 881 => bit_in_tb <= '1';
                WHEN 882 => bit_in_tb <= '1';
                WHEN 883 => bit_in_tb <= '0';
                WHEN 884 => bit_in_tb <= '0';
                WHEN 885 => bit_in_tb <= '1';
                WHEN 886 => bit_in_tb <= '0';
                WHEN 887 => bit_in_tb <= '1';
                WHEN 888 => bit_in_tb <= '0';
                WHEN 889 => bit_in_tb <= '1';
                WHEN 890 => bit_in_tb <= '1';
                WHEN 891 => bit_in_tb <= '0';
                WHEN 892 => bit_in_tb <= '1';
                WHEN 893 => bit_in_tb <= '0';
                WHEN 894 => bit_in_tb <= '1';
                WHEN 895 => bit_in_tb <= '0';
                WHEN 896 => bit_in_tb <= '0';
                WHEN 897 => bit_in_tb <= '1';
                WHEN 898 => bit_in_tb <= '1';
                WHEN 899 => bit_in_tb <= '0';
                WHEN 900 => bit_in_tb <= '0';
                WHEN 901 => bit_in_tb <= '1';
                WHEN 902 => bit_in_tb <= '1';
                WHEN 903 => bit_in_tb <= '0';
                WHEN 904 => bit_in_tb <= '1';
                WHEN 905 => bit_in_tb <= '1';
                WHEN 906 => bit_in_tb <= '1';
                WHEN 907 => bit_in_tb <= '0';
                WHEN 908 => bit_in_tb <= '1';
                WHEN 909 => bit_in_tb <= '0';
                WHEN 910 => bit_in_tb <= '1';
                WHEN 911 => bit_in_tb <= '0';
                WHEN 912 => bit_in_tb <= '1';
                WHEN 913 => bit_in_tb <= '0';
                WHEN 914 => bit_in_tb <= '0';
                WHEN 915 => bit_in_tb <= '0';
                WHEN 916 => bit_in_tb <= '0';
                WHEN 917 => bit_in_tb <= '1';
                WHEN 918 => bit_in_tb <= '0';
                WHEN 919 => bit_in_tb <= '0';
                WHEN 920 => bit_in_tb <= '0';
                WHEN 921 => bit_in_tb <= '0';
                WHEN 922 => bit_in_tb <= '1';
                WHEN 923 => bit_in_tb <= '0';
                WHEN 924 => bit_in_tb <= '0';
                WHEN 925 => bit_in_tb <= '1';
                WHEN 926 => bit_in_tb <= '1';
                WHEN 927 => bit_in_tb <= '1';
                WHEN 928 => bit_in_tb <= '0';
                WHEN 929 => bit_in_tb <= '0';
                WHEN 930 => bit_in_tb <= '1';
                WHEN 931 => bit_in_tb <= '0';
                WHEN 932 => bit_in_tb <= '1';
                WHEN 933 => bit_in_tb <= '1';
                WHEN 934 => bit_in_tb <= '0';
                WHEN 935 => bit_in_tb <= '1';
                WHEN 936 => bit_in_tb <= '1';
                WHEN 937 => bit_in_tb <= '0';
                WHEN 938 => bit_in_tb <= '1';
                WHEN 939 => bit_in_tb <= '0';
                WHEN 940 => bit_in_tb <= '1';
                WHEN 941 => bit_in_tb <= '0';
                WHEN 942 => bit_in_tb <= '1';
                WHEN 943 => bit_in_tb <= '0';
                WHEN 944 => bit_in_tb <= '1';
                WHEN 945 => bit_in_tb <= '1';
                WHEN 946 => bit_in_tb <= '1';
                WHEN 947 => bit_in_tb <= '0';
                WHEN 948 => bit_in_tb <= '1';
                WHEN 949 => bit_in_tb <= '1';
                WHEN 950 => bit_in_tb <= '0';
                WHEN 951 => bit_in_tb <= '1';
                WHEN 952 => bit_in_tb <= '1';
                WHEN 953 => bit_in_tb <= '0';
                WHEN 954 => bit_in_tb <= '0';
                WHEN 955 => bit_in_tb <= '0';
                WHEN 956 => bit_in_tb <= '1';
                WHEN 957 => bit_in_tb <= '0';
                WHEN 958 => bit_in_tb <= '0';
                WHEN 959 => bit_in_tb <= '0';
                WHEN 960 => bit_in_tb <= '1';
                WHEN 961 => bit_in_tb <= '1';
                WHEN 962 => bit_in_tb <= '0';
                WHEN 963 => bit_in_tb <= '1';
                WHEN 964 => bit_in_tb <= '1';
                WHEN 965 => bit_in_tb <= '0';
                WHEN 966 => bit_in_tb <= '1';
                WHEN 967 => bit_in_tb <= '0';
                WHEN 968 => bit_in_tb <= '1';
                WHEN 969 => bit_in_tb <= '1';
                WHEN 970 => bit_in_tb <= '1';
                WHEN 971 => bit_in_tb <= '1';
                WHEN 972 => bit_in_tb <= '0';
                WHEN 973 => bit_in_tb <= '1';
                WHEN 974 => bit_in_tb <= '1';
                WHEN 975 => bit_in_tb <= '1';
                WHEN 976 => bit_in_tb <= '1';
                WHEN 977 => bit_in_tb <= '1';
                WHEN 978 => bit_in_tb <= '0';
                WHEN 979 => bit_in_tb <= '0';
                WHEN 980 => bit_in_tb <= '1';
                WHEN 981 => bit_in_tb <= '1';
                WHEN 982 => bit_in_tb <= '1';
                WHEN 983 => bit_in_tb <= '0';
                WHEN 984 => bit_in_tb <= '1';
                WHEN 985 => bit_in_tb <= '1';
                WHEN 986 => bit_in_tb <= '0';
                WHEN 987 => bit_in_tb <= '0';
                WHEN 988 => bit_in_tb <= '0';
                WHEN 989 => bit_in_tb <= '0';
                WHEN 990 => bit_in_tb <= '0';
                WHEN 991 => bit_in_tb <= '1';
                WHEN 992 => bit_in_tb <= '0';
                WHEN 993 => bit_in_tb <= '0';
                WHEN 994 => bit_in_tb <= '0';
                WHEN 995 => bit_in_tb <= '1';
                WHEN 996 => bit_in_tb <= '0';
                WHEN 997 => bit_in_tb <= '1';
                WHEN 998 => bit_in_tb <= '1';
                WHEN 999 => bit_in_tb <= '1';
                WHEN 1000 => bit_in_tb <= '0';
                WHEN 1001 => bit_in_tb <= '0';
                WHEN 1002 => bit_in_tb <= '0';
                WHEN 1003 => bit_in_tb <= '0';
                WHEN 1004 => bit_in_tb <= '0';
                WHEN 1005 => bit_in_tb <= '1';
                WHEN 1006 => bit_in_tb <= '1';
                WHEN 1007 => bit_in_tb <= '0';
                WHEN 1008 => bit_in_tb <= '1';
                WHEN 1009 => bit_in_tb <= '1';
                WHEN 1010 => bit_in_tb <= '0';
                WHEN 1011 => bit_in_tb <= '1';
                WHEN 1012 => bit_in_tb <= '1';
                WHEN 1013 => bit_in_tb <= '1';
                WHEN 1014 => bit_in_tb <= '0';
                WHEN 1015 => bit_in_tb <= '0';
                WHEN 1016 => bit_in_tb <= '1';
                WHEN 1017 => bit_in_tb <= '0';
                WHEN 1018 => bit_in_tb <= '0';
                WHEN 1019 => bit_in_tb <= '1';
                WHEN 1020 => bit_in_tb <= '0';
                WHEN 1021 => bit_in_tb <= '0';
                WHEN 1022 => bit_in_tb <= '1';
                WHEN 1023 => bit_in_tb <= '0';
               WHEN	OTHERS	=>	NULL;
           END CASE;
           if count >= 1024 then
               bit_in_tb <= 'Z';
           end if;
           if count = len then testing <= false;      -- fine test
           end if;
           if (count >= len) then NULL;
           end if;
           count <= count + 1;
       end if;


end process proc_test;

end interleaver_test;
